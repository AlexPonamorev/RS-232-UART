	/* имеем данные на шине приема передающиеся с частотой 115200 - заранее декларированной.
	 имеем опороную частоту тактирование схемы clk_i == 50_000_000 Гц - CLK_FREQ
	 для приема данных необходим счетчик считающий до Cout_Clk == CLK_FREQ/ 115200 в интервале счета от cntrl== 0  до значения  &cntrl == 1 - имеем период принимаемого бита как Counter_Div_Clk_Rx == Cout_Clk
	 принимаемые данные перенесены в клоковый домен приемника регистром Reg_Synchron на выходе которого имеем данные - готовые для обработки приемником. 
	 создадим счетчик длины принимаемого бита Counter_Int_Bit - для записи выборки с шины в регистр сдвига для дальнейшего анализа в мажоритарной схеме
	 за такт до такта коэффициента деления анализируем мажоритарную схему и определяем флаг записи start
	 запись в сдвиговый регистр на средине принимаемого бита
	*/
module Uart_RX_1318
	
 (
	// control
	input            Clk_RX ,                           // тактовый сигнал приемника 50_000_000
	input            Reset_R ,
	// RS-232 interface
	input            DATA_RX_In ,                        //входная несинхронизированная шина данных
	// user signals
	output reg     Ok_Data_Rx                           // сигнал готовности для считывания принятого байта с регистра
	output[7:0]    DATA_RX_Out              
);
	localparam Cout_Clk  = (CLK_FREQ / BAUD_RATE);       // значение, по достижению котогого счетчиком делителя -выдаем управляющий сигнал на схему 
    localparam Cout_Bit = clob2(Cout_Clk);               //параметр для вычисления разрядности счетчика делителя частот
	
	parameter BAUD_RATE  = 115200;
	parameter CLK_FREQ   = 50_000_000;
	parameter Parity_Bit = 1'b1;
	parameter Stop_Bit   = 1'b1;
	
	reg  [3:0] Counter_Rec_Bit;                          // счетчик принятых бит -разрядность беру с запасом для дальнейшей доработки
	reg  [2:0] Reg_Synchron;                   			 // регистр переноса данных в в клоковый домен модуля 
	wire       RX_Synchron;                         	 //синхронизированная с частотой модуля линия данных
	
	reg  [2:0] Shift_Maj;                                //сдвиговый регистр выборки данных
	reg  [1:0] Counter_Int_Bit;                          //счетчик битовых интервалов (кол-ва периодов)
	wire       Maj_Data ;                                // валидности нуля на шине
	reg        start;                                    // регистр хранения результата проверки линни на старт бит
	reg        Xor_Valid;                                // регистр хранения результата проверки на четность
	reg        Stop_Bit_Valid;                           // регистр хранения результата проверки на Stop_Bit
	
	reg [7 + Stop_Bit + Parity_Bit:0] R_Shift_DATA_RX;  // регистр для приема байта 
/**********************************************************************************************************************/
	//несентизируемый блок,функция вычисления разрядности счетчика делителя частот// количество D триггеров // разрядность - функция log2 чтобы получить нужное кол-во триггеров для счета
	function integer clob2(input[31:0] value );
		if (value < 2)
		clob2 = 1;
	else 
		begin
			value = value - 1;
			for (clob2 = 0; value > 0; clob2 = clob2 + 1)
			value = value >> 1;      
		end
	endfunction
	
	reg [Cout_Bit-1:0] Counter_Div_Clk_Rx;  // счетчик делитель частот  
/**********************************************************************************************************************/
	// модуль для синхронизации входной частоты приема        
	always @(posedge Clk_RX)	
	begin
		if(~Reset_R)
		Reg_Synchron <= {3{1'b1}};  //состояние готовности к работе
		else                                                             // И НА ТАКТЕ КОЭФФ ДЕЛЕНИЯ
		Reg_Synchron <= {DATA_RX_In,Reg_Synchron[2:1]};              //со младшего выдаем
	end
	
	assign RX_Synchron = Reg_Synchron[0];
/*****************************************************************************************************************************/
	// счетчик инкрементируется до значения == коэффициенту от деления частот являимущяся ТАКТОМ для работы схемы ,  обеспечивающим нужную частоту приема - Counter_Div_Clk_Rx == Cout_Clk 115200
	//счетчик делитель частот           
	always@(posedge Clk_RX)
	begin
		if (~Reset_R || Counter_Div_Clk_Rx == Cout_Clk)
		Counter_Div_Clk_Rx <= {(Cout_Bit-1){1'b0}};          //скинуть счетчик в нуль                                 
		else
		Counter_Div_Clk_Rx <= Counter_Div_Clk_Rx + 1'b1 ;                                          
	end
/********************************************************************************************************************************************************************************************/
	//счетчик делитель принимаемого бита
	//счетчик инкрементируется cntr + 1 на частоте деления  Cout_Clk/3   
	always@(posedge Clk_RX)
		if (~Reset_R || (RX_Synchron == 1'b0 && Counter_Rec_Bit == 4'b1111) || Counter_Int_Bit == 2'd2) // после инициализации и последущей проверки на данные условия постоянно сбрасывается в  4'b000  
		Counter_Int_Bit <= 2'b0;
		else if  (Counter_Div_Clk_Rx == Cout_Clk-1/3)           
		Counter_Int_Bit <= Counter_Int_Bit + 1'b1;
/********************************************************************************************************************************************************************************************/
	//счетчик принятых бит //на восьмом такте ожидаем Stop_Bit 
	always@(posedge Clk_RX)
		if (~Reset_R || (Counter_Rec_Bit == (4'd8 + Stop_Bit + Parity_Bit) && Counter_Div_Clk_Rx == Cout_Clk))  // последнее условие - переход в режим ожидания - т.е позицию старта 
			Counter_Rec_Bit <= 4'b1111;                        //стартовая позиция
		else if (start == 1'b0 && Counter_Div_Clk_Rx == Cout_Clk - 1 )     
		    Counter_Rec_Bit <= Counter_Rec_Bit + 1'b1;
/*********************************************************************************************************************************************************************************************/
	//мажоритарноя выборка - схема определяющая начало приема // работае от счетчика интервалов
	always@(posedge Clk_RX)   
		if (~Reset_R && Counter_Rec_Bit == (4'd8 + Stop_Bit + Parity_Bit))
			Shift_Maj <= {3{1'b1}};   
		else if(Counter_Int_Bit == 2'd0 || Counter_Int_Bit == 2'd1 || Counter_Int_Bit == 2'd2)  // задвигаем в регистр для  мажоритарного анализа того что приняли
		   Shift_Maj <= {RX_Synchron,Shift_Maj[2:1]};
	 
	assign Maj_Data = Shift_Maj[0] & Shift_Maj[1] | Shift_Maj[0] | Shift_Maj[2] |Shift_Maj[1] & Shift_Maj[2]; //анализ принятого бита
/***********************************************************************************************************************************************************************************************/
	//флаг валидности нуля шины   -  старт отсчета для счетчика принятых бит 	   
	always@(posedge Clk_RX)
			if(~Reset_R && Counter_Rec_Bit == 4'b1111)
			start <= 1'b1;
			else if (Maj_Data == 1'b0 && Counter_Div_Clk_Rx == Cout_Clk - 1'b1) //  за один такт до обнуления счетчика интервалов, так как со следующего такта нужно уже иметь какое то значение на регистре старта
			start <= 1'b0;
/************************************************************************************************************************************************************************************************/		
	// регистр принимаемого байта
	always@(posedge Clk_RX)
		if (~Reset_R)
		R_Shift_DATA_RX <= {(8 + Stop_Bit + Parity_Bit){1'b1}};
		else if (start == 1'b0 && Counter_Int_Bit == 2'd1 && Counter_Rec_Bit < 4'd9 + Stop_Bit + Parity_Bit )  // на середине бита записать значение на шине
		
		R_Shift_DATA_RX <= {RX_Synchron,R_Shift_DATA_RX[7 + Parity_Bit + Stop_Bit:1]};
/*************************************************************************************************************************************************************************************************/
	// вычисление валидности принятого байта 
	always@(posedge Clk_RX)
		if (~Reset_R || Counter_Rec_Bit == 4'b1111)
		Ok_Data_Rx <= 1'b0;                          // в состоянии отсутствия данных 
	else if (Counter_Rec_Bit == 4'd8 + Stop_Bit + Parity_Bit && Counter_Div_Clk_Rx == Cout_Clk-1 && Maj_Data == 1'b1 && Xor_Valid == 1'b1 && Stop_Bit_Valid == 1'b1)
		begin
			Ok_Data_Rx <= 1'b1;                          // разрешение на считывание из байта 
			start <= 1'b0;                                // вернем старт в режим ожидания
		end
		
	assign DATA_RX_Out[7:0]= R_Shift_DATA_RX[7:0];              
	assign Xor_Data_RX = ^R_Shift_DATA_RX[7:0];
	
/****************************************************************************************************************************************/
//                              костыль для реализации проверки на четность
//на восьмом такте имеем некое значение функции четности по регистру [7:0] в котором находится байт данных
//на этом же такте сравниваем значение в восьмом регистре байта с вычисленным значение по [7:0] 
//на девятом такте (по факту он десятый т.к.отчсчет с нуля) в зависимости от предыдущего результа записываем "0" либо "1" в регистр хранениячетности
	always@(posedge Clk_RX)
	begin
		if(~Reset_R || Counter_Rec_Bit == 4'b1111 )
		Xor_Valid <= 1'b0;
		else if(Parity_Bit == 1'b1 && Counter_Rec_Bit == 4'd8 &&  Counter_Div_Clk_Rx == Cout_Clk - 1)
			begin
				if((R_Shift_DATA_RX[8] == Xor_Data_RX)
				Xor_Valid <= 1'b1;
				else
				Xor_Valid <= 1'b0;
			end	   
		else
	    Xor_Valid <= 1'b1;                          // во всех остальных случаях будем считать что он есть
		   
	end	
	
/***********************************************************************************************************************************************************/
//      					   повторяю описанный ранее алгоритм в отношении стоп бита
	 always@(posedge Clk_RX)
	begin
		if(~Reset_R ||Counter_Rec_Bit == 4'b1111 )
		Stop_Bit_Valid <= 1'b0;
		else if(Stop_Bit == 1'b1 && Counter_Rec_Bit == 4'd8 &&  Counter_Div_Clk_Rx == Cout_Clk - 1)
			begin
				if((R_Shift_DATA_RX[9] == Xor_Data_RX)
				Stop_Bit_Valid <= 1'b1;
				else
				Stop_Bit_Valid <= 1'b0;                  
			end	   
		else
	    Stop_Bit_Valid <= 1'b1;                         // во всех остальных случаях будем считать что он есть   
		   
	end	




	
	















endmodule