module Uart_TX_1318( 
	input Clk_TX ,                                   // опорная частота                                    
	input Reset_T,                                   // сброс,активен по "0" 
	input Start,                                     // линия сигнала на  записи байта в передатчик (внешний старт передатчика)
	input [7:0] Data_TX_In,                          // восьмибитный вход на приемник
	output Ena_New_Data,                             // флаг состояния готовности к работе
	output TX_Out                                    // последовательный выход на передатчик
	);
	
	parameter CLK_FREQ_T  = 100_000_000;              // входная частота          // параметр внешний                               
	parameter BAUD_RATE   = 115200;                   // желаемая частота передачи пакета  // параметр внешний                   
	parameter Parity_Bit  = 1'b1;                     // наличие бита четности( либо есть ,либо нет -> 1'b1 || 1'b0 )
	parameter Stop_Bit    = 1'b1;                     // наличие и длинна стоп бита       
	localparam Cout_Clk_T = CLK_FREQ_T/BAUD_RATE;     // коэфициент деления частот        
	localparam Cout_Bit_T = Clob2(Cout_Clk_T);        // параметр для вычисления разрядности счетчика делителя частот       


	reg [3:0] Count_Bit;                              //регистр счетчика выгрузки пакета             
	reg [8 + Parity_Bit:0] Reg_Shift_Data;            // регистр пакета данных         
	reg [Cout_Bit_T-1:0]  Counter_Div_clk;            // регистр счетчика делителя частот     
	wire Start_Front;                                 // внутренний старт формируется по перепаду внешнего с 0 в 1 
	reg Reg_Srart_Front ;                             // регистр для формирования фронта внутреннего старта
	wire Start_0;                                     // техническое соединение
	wire Xor_Data_TX;                                 // элемент для вычисления четности в пакете данных                              
	 
	//******************************************************************************************** //
	//несентизируемый блок,функция вычисления разрядности счетчика делителя частот// количество D триггеров //как функция log2(по основанию 2)
	function integer Clob2(input[31:0] value );
		if (value < 2)
		Clob2 = 1;
	else 
		begin
		value = value - 1;
		for (Clob2 = 0; value > 0; Clob2 = Clob2 + 1)
		value = value >> 1;      
		end
	endfunction



//***************************************************************************************************//
//  счетчик делитель частот
	always @ (posedge  Clk_TX) 
		if (~Reset_T || Counter_Div_clk == Cout_Clk_T || Start_Front )          // Counter_Div_clk == Cout_Clk_T//значение счетчика равна коэфф. деления                 
		Counter_Div_clk <= {(Count_Bit-1) {1'b0}};                            // обеспечивает выдачу бита с региста каждые 115200 тактов                                         
	else
		Counter_Div_clk <= Counter_Div_clk + 1'b1 ;                                  
 

//***************************************************************************************************//
//тело регистра пакета данных (ТЛПД) структура- линия передачи в отсутствии данных всегда в ...1'b1...(вседа выгружается)/стоп бит(1)/бит четности/пакет данных/старт бит (всегда 1'b0)/в 1'b1...
	always @(posedge  Clk_TX)               //    стоп бит и его длинна определяется работой СВ !!!                                     ->ст.регистр->>>>>>>>>>>>>>>>>>>>>>>>>мл.рег.->
		begin
		if (~Reset_T)
		Reg_Shift_Data <= {8 + Parity_Bit{1'b1}};                                  //записать ТЛПД единицы // в 8 регистров + регистр бита четности ->положить единицы                           
	else if (Start_Front)                                                            // по внутреннему старту - т.к. он будет всегда  длительностью в clock  вне зависимости от длительности внешнего старта                    
		Reg_Shift_Data <= {(Parity_Bit ? Xor_Data_TX : 1'b1) , Data_TX_In, 1'b0};              // в зависимотсти от наличия бита четности в старший разряд регистра будет положено либо значение функции четности                    
	else if(Counter_Div_clk == Cout_Clk_T && Count_Bit < 4'h9 + Stop_Bit + Parity_Bit ) //либо единица, которая также может быть стоп битом        
		 Reg_Shift_Data <=  {1'b1 , Reg_Shift_Data[8 + Parity_Bit :1]};              // в старший разряд заполнить 1'b1             
	end
  
	assign TX_Out = Reg_Shift_Data[0];
 //*****************************************************************************************************//
 // счетчик выгрузки ТЛПД (СВ)
	always @ (posedge  Clk_TX)
		 if(~Reset_T ) 
		Count_Bit <= 4'h9 + Parity_Bit + Stop_Bit;                               // счетчик по умолчанию хранит это значение 
	else if ( Start_Front && Ena_New_Data )                                                    // по сигналу внутреннего старта и разрешения сбрасывается в нуль
		Count_Bit <= 1'b0;
	else if (Counter_Div_clk == Cout_Clk_T && Count_Bit < 4'h9 + Stop_Bit + Parity_Bit) // инкрементировать счетчик пока счетчик делителя не дойдет до значения коэфициента деления и(&&)
                                                                                  //и счетчик выгрузки не дойдет до требуемого значения( в зависимости от параметров)                                                                                                                                                                 
                     Count_Bit <=Count_Bit + 1'b1;                                   
                                                                                                                      
	else if (Count_Bit == 4'h9 && Counter_Div_clk == Cout_Clk_T && (Parity_Bit || Stop_Bit))         
		Count_Bit <= (4'h9 + Parity_Bit + Stop_Bit);
	else 
		Count_Bit <= Count_Bit; 

 //*******************************************************************************************************//
 //блок генерации сигнала разрешения 

	assign Ena_New_Data = !(Count_Bit < 4'h9 + Stop_Bit + Parity_Bit);

//*********************************************************************************************************//
//блок генерации фронта внутреннего старта // защита от залипания внешнего старта
	always @(posedge  Clk_TX )
		begin
		if (~Reset_T  )
		Reg_Srart_Front <= 0;              
	else         
		Reg_Srart_Front <= Start_0;                                  
		end
		
	assign Start_0 = Ena_New_Data ? Start : 1'b0 ;     //защита от подачи старта     
	assign Start_Front = ~Reg_Srart_Front & Start_0;   //выделяем фронт
//************************************************************************************************************//
// реализация вычисления четности байта(регистра)	
		assign Xor_Data_TX = ^ Data_TX_In ;                   

endmodule 